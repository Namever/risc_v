module DE0_CV(

	//////////// CLOCK //////////
	input 		          		CLOCK_50,
	input 		          		CLOCK2_50,
	input 		          		CLOCK3_50,
	inout 		          		CLOCK4_50,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,

	//////////// SEG7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
	output		     [6:0]		HEX2,
	output		     [6:0]		HEX3,
	output		     [6:0]		HEX4,
	output		     [6:0]		HEX5,

	//////////// KEY //////////
	input 		     [3:0]		KEY,
	input 		          		RESET_N,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// PS2 //////////
	inout 		          		PS2_CLK,
	inout 		          		PS2_CLK2,
	inout 		          		PS2_DAT,
	inout 		          		PS2_DAT2,

	//////////// microSD Card //////////
	output		          		SD_CLK,
	inout 		          		SD_CMD,
	inout 		     [3:0]		SD_DATA,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// VGA //////////
	output		     [3:0]		VGA_B,
	output		     [3:0]		VGA_G,
	output		          		VGA_HS,
	output		     [3:0]		VGA_R,
	output		          		VGA_VS,

	//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
	inout 		    [35:0]		GPIO_0,

	//////////// GPIO_1, GPIO_1 connect to GPIO Default //////////
	inout 		    [35:0]		GPIO_1
);

//=======================================================
//  REG/WIRE declarations
//=======================================================


//`define Burn
logic [31:0] regs_31;
logic clk;
logic clk_div;

//=======================================================
//  Structural coding
//=======================================================
`ifdef Burn

clock_divider u_clock_divider(
    .clk    (CLOCK_50),
    .rst    (~RESET_N),
    .DIVISOR(10000),
    .clk_out(clk_div)
);

assign clk = clk_div;
`else
assign clk = CLOCK_50;
`endif

Top u_Core(
    .clk    (clk),
    .rst    (~RESET_N),
    .regs_31(regs_31)
);

// Instance for 7-segment display for each HEX display
seven_segment_display u_seven_0(
	.digit (regs_31[3:0]),
	.seg (HEX0)
);

seven_segment_display u_seven_1(
	.digit (regs_31[7:4]),
	.seg (HEX1)
);

seven_segment_display u_seven_2(
	.digit (regs_31[11:8]),
	.seg (HEX2)
);

seven_segment_display u_seven_3(
	.digit (regs_31[15:12]),
	.seg (HEX3)
);

seven_segment_display u_seven_4(
	.digit (regs_31[19:16]),
	.seg (HEX4)
);

seven_segment_display u_seven_5(
	.digit (regs_31[23:20]),
	.seg (HEX5)
);


// Assign `regs_31`[9:0] to LEDs
assign LEDR = regs_31[9:0];

endmodule
